module pri_en83_tb();
reg[7:0] a;
wire[2:0] y;
pri_en83 i1(a,y);
initial 
begin
        a=8'b0000_0000;
    #10 a=8'b0000_0001;
    #10 a=8'b0000_0010;
    #10 a=8'b0000_0101;
    #10 a=8'b0000_1001;
    #10 a=8'b0001_0010;
    #10 a=8'b0010_0000;
    #10 a=8'b0100_1100;
    #10 a=8'b1000_0000;
end
endmodule
